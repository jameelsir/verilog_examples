`timescale 1ns / 1ps

module tb_mux2x1;

    // Inputs
    reg a;
    reg b;
    reg sel;

    // Output
    wire y;

    // Instantiate the Unit Under Test (UUT)
    mux2x1 uut (
        .a(a),
        .b(b),
        .sel(sel),
        .y(y)
    );

    initial begin
        // Initialize waveform dump
        $dumpfile("tb_mux2x1.vcd");
        $dumpvars(0, tb_mux2x1);

        // Initialize Inputs
        a = 0; b = 0; sel = 0;

        // Test all input combinations
        #10 a = 0; b = 0; sel = 0;
        #10 a = 0; b = 1; sel = 0;
        #10 a = 1; b = 0; sel = 0;
        #10 a = 1; b = 1; sel = 0;
        #10 a = 0; b = 0; sel = 1;
        #10 a = 0; b = 1; sel = 1;
        #10 a = 1; b = 0; sel = 1;
        #10 a = 1; b = 1; sel = 1;
        #10;

        $finish;
    end

    initial begin
        $monitor("Time=%0t | a=%b b=%b sel=%b | y=%b", $time, a, b, sel, y);
    end

endmodule